module alu_ctrl (
    input  logic [2:0] funct3_i,
    input  logic [6:0] funct7_i,
    input  logic [1:0] alu_ctrl_i,
    output logic [3:0] alu_op_o
);

endmodule
