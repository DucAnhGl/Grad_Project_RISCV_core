module insn_vld_dec (
    input  logic [31:0] instr_i,
    output logic insn_vld_o
);



endmodule